`timescale 1ns / 1ps
module shifteru0(
	input [47:0] u0,
	input [5:0] exp_e,
	output reg [47:0] x_e
);

always @(exp_e or u0) begin
case(exp_e)
	1: x_e <= u0 << 1;
	2: x_e <= u0 << 2;
	3: x_e <= u0 << 3;
	4: x_e <= u0 << 4;
	5: x_e <= u0 << 5;
	6: x_e <= u0 << 6;
	7: x_e <= u0 << 7;
	8: x_e <= u0 << 8;
	9: x_e <= u0 << 9;
	10: x_e <= u0 << 10;
	11: x_e <= u0 << 11;
	12: x_e <= u0 << 12;
	13: x_e <= u0 << 13;
	14: x_e <= u0 << 14;
	15: x_e <= u0 << 15;
	16: x_e <= u0 << 16;
	17: x_e <= u0 << 17;
	18: x_e <= u0 << 18;
	19: x_e <= u0 << 19;
	20: x_e <= u0 << 20;
	21: x_e <= u0 << 21;
	22: x_e <= u0 << 22;
	23: x_e <= u0 << 23;
	24: x_e <= u0 << 24;
	25: x_e <= u0 << 25;
	26: x_e <= u0 << 26;
	27: x_e <= u0 << 27;
	28: x_e <= u0 << 28;
	29: x_e <= u0 << 29;
	30: x_e <= u0 << 30;
	31: x_e <= u0 << 31;
	32: x_e <= u0 << 32;
	33: x_e <= u0 << 33;
	34: x_e <= u0 << 34;
	35: x_e <= u0 << 35;
	36: x_e <= u0 << 36;
	37: x_e <= u0 << 37;
	38: x_e <= u0 << 38;
	39: x_e <= u0 << 39;
	40: x_e <= u0 << 40;
	41: x_e <= u0 << 41;
	42: x_e <= u0 << 42;
	43: x_e <= u0 << 43;
	44: x_e <= u0 << 44;
	45: x_e <= u0 << 45;
	46: x_e <= u0 << 46;
	47: x_e <= u0 << 47;
	48: x_e <= u0 << 48;
	default: x_e <= u0;
endcase
end
endmodule
	

