`timescale 1ns / 1ps
module shiftere(
	input [30:0] e,
	input [5:0] exp_f,
	output reg [30:0] x_f1 
);

always @(exp_f or e) begin
case(exp_f)
	6'b000101: x_f1 <= e >> 5;
	6'b000100: x_f1 <= e >> 4;
	6'b000011: x_f1 <= e >> 3;
	6'b000010: x_f1 <= e >> 2;
	6'b000001: x_f1 <= e >> 1;
	6'b000000: x_f1 <= e;
	6'b111111: x_f1 <= e << 1;
	6'b111110: x_f1 <= e << 2;
	6'b111101: x_f1 <= e << 3;
	6'b111100: x_f1 <= e << 4;
	6'b111011: x_f1 <= e << 5;
	6'b111010: x_f1 <= e << 6;
	6'b111001: x_f1 <= e << 7;
	6'b111000: x_f1 <= e << 8;
	6'b110111: x_f1 <= e << 9;
	6'b110110: x_f1 <= e << 10;
	6'b110101: x_f1 <= e << 11;
	6'b110100: x_f1 <= e << 12;
	6'b110011: x_f1 <= e << 13;
	6'b110010: x_f1 <= e << 14;
	6'b110001: x_f1 <= e << 15;
	6'b110000: x_f1 <= e << 16;
	6'b101111: x_f1 <= e << 17;
	6'b101110: x_f1 <= e << 18;
	6'b101101: x_f1 <= e << 19;
	6'b101100: x_f1 <= e << 20;
	6'b101011: x_f1 <= e << 21;
	6'b101010: x_f1 <= e << 22;
	6'b101001: x_f1 <= e << 23;
	6'b101000: x_f1 <= e << 24;
	6'b100111: x_f1 <= e << 25;
	default: x_f1 <= e;
endcase
end

endmodule
